.MODEL BC547C NPN( 
+     IS=4.679E-14
+     NF=1.01
+     ISE=2.642E-15
+     NE=1.581
+     BF=458.7
+     IKF=0.1371
+     VAF=52.64
+     NR=1.019
+     ISC=2.337E-14
+     NC=1.164
+     BR=11.57
+     IKR=0.1144
+     VAR=364.5
+     RB=1
+     IRB=1E-06
+     RBM=1
+     RE=0.2598
+     RC=1
+     XTB=0
+     EG=1.11
+     XTI=3
+     CJE=1.229E-11
+     VJE=0.5591
+     MJE=0.3385
+     TF=4.689E-10
+     XTF=160
+     VTF=2.828
+     ITF=0.8842
+     PTF=0
+     CJC=4.42E-12
+     VJC=0.1994
+     MJC=0.2782
+     XCJC=0.6193
+     TR=1E-32
+     CJS=0
+     VJS=0.75
+     MJS=0.333
+     FC=0.7936 )
*
