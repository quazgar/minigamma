* (vin)----R1---(1)---R2----(-)

Vin vin 0 pulse 9 0.6 1u 100n 100n 1u
R1 vin 1 100k
R2 1 0 200k
  
.end
