* (vin)----R1(1000)---(1)   //// ---R2(100)----(-)
*                     |
*                    C1(1uF)----------(-)
*
* => tau = 1ms

Vin vin 0 pulse 0 1 0.2u 100n 100n 1.5m
R1 vin 1 1000
*R2 1 0 100
C1 1 0 1u

.end
