.MODEL BC557 PNP(
* + IS=3.834E-14
* + NF=1.008
* + ISE=1.219E-14
* + NE=1.528
* + BF=800
* + IKF=0.08039
* + VAF=21.11
* + NR=1.005
* + ISC=2.852E-13
* + NC=1.28
* + BR=14.84
* + IKR=0.047
* + VAR=32.02
* + RB=1
* + IRB=1E-06
* + RBM=1
* + RE=0.6202
* + RC=0.5713
* + XTB=0
* + EG=1.11
* + XTI=3
* + CJE=1.23E-11
* + VJE=0.6106
* + MJE=0.378
* + TF=5.595E-10
* + XTF=3.414
* + VTF=5.23
* + ITF=0.1483
* + PTF=0
* + CJC=1.084E-11
* + VJC=0.1022
* + MJC=0.3563
* + XCJC=0.6288
* + TR=1E-32
* + CJS=0
* + VJS=0.75
* + MJS=0.333
* + FC=0.8027 )
+ BF=800
+)
